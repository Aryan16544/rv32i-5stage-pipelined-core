`timescale 1ns / 1ps

module register_file (
    input  wire        clk,
    input  wire        rst,

    input  wire [4:0]  rs1,
    input  wire [4:0]  rs2,

    input  wire [4:0]  rd,
    input  wire        rd_we,
    input  wire [31:0] rd_data,

    output wire [31:0] rs1_data,
    output wire [31:0] rs2_data
);

    reg [31:0] regs [0:31];
    integer i;

    // Reset
    always @(posedge clk) begin
        if (rst) begin
            for (i = 0; i < 32; i = i + 1)
                regs[i] <= 32'b0;
        end else if (rd_we && rd != 5'd0) begin
            regs[rd] <= rd_data;
        end
    end

    assign rs1_data = (rs1 == 5'd0) ? 32'b0 : regs[rs1];
    assign rs2_data = (rs2 == 5'd0) ? 32'b0 : regs[rs2];

endmodule
